-------------------------------------------------------------------------------
-- (start) add2_flat_tb.vhd
-------------------------------------------------------------------------------
-- Question 8

library ieee;
use ieee.std_logic_1164.all;

  -- insert VHDL testbench code here


-- Question 8(c)
  --insert answer here

-- Question 8(e)
  --insert answer here

-------------------------------------------------------------------------------
-- (end) add2_flat_tb.vhd
-------------------------------------------------------------------------------
